ifndefGUARDAMBA DEFS SVHdefineGUARD AMBA DEFS SVH
defineDC SRESP WDdefine RESP ERRBUS WDdefine SLV CFG ADDR WD
23
// AHB/AXI response data width// The width of encoded error response bus
32
// programmable width used to select the address range for
confiquration
define SLV IO ADDR WD
// programmable width used to select the address range for IO
32
transaction
define MSTR CFG ADDR WD
// programmable width used to select the address range for
32
configuration
define MSTR IO ADDR WD
32
// programmable width used to select the address range for IO
transaction
// 5bits type， 3bits TC， 2bits Attr， 5 bits IO,ROMand MEMBAR//define MSTR MISC INFO WD(5+3+2+5+3+3+3)range, 3bits function number, 3bits of status, 3bits of byte length offsetdefine MSTR MISC INFO TYPE HIGH
23191816151413106532e
define MSTR MISC INFO TYPE LOWdefine MSTR MISC INFO TC HIGHdefine MSTR MISC INFO TC LOWdefine MSTR MISC INFO ATTR HIGHdefine MSTR MISC INFO ATTR LOWdefineMSTR MISC INFO FUNC HIGH
define MSTR MISC INFO FUNC LOWdefine MSTR MISC INFO BAR HIGH
define MSTR MISC INFO BAR LOWdefine MSTR MISC INFO STATUS HIGH
define MSTR MISC INFO STATUS LOWdefine MSTR MISC INFO LEN OFFSET HIGHdefine MSTR MISC INFO LEN OFFSET LOW
define MSTR MISC INFO REOID LOWdefine MSTR MISC INFO REQID HIGHdefine MSTR MISC INFO TAG LOW
define MSTR MISC INFO TAG HIGH
MSTR MISC INFO TYPE HIGH + 1MSTR MISC INFO REQID LOW +16“MSTR MISC INFO REQID HIGH + 1MSTR MISC INFO TAG LOW +8- 1
define MSTR MISC INFO VF HIGHMSTR MISC INFO TAG HIGHMSTR MISC INFO VF HIGHdefine MSTR MISC INFO ATS NWMSTR MISC INFO PE HIGH/'define SLV RESP MISC INFO WD(1+3+3+2+1+1+3)2bits Attr. l bit TD and 1 Bit BCM 3 Bit Func Num
define MSTR MISC INFO PF HIGH
// lbit for response of NP write, 3bits status, 3bits TC,
-------------
---------
associate to SLV MISC INFO WD
----------- NOte ---------------------The SLV MISC INFO WD has been moved to AMBA cc constant because of a script issue/ please update the amba cc constant file in future when this busgrows/ifdef AHB POPULATED/define SLV MISC INFO WD(1+ 4 + 8 + 3 + 2 +1+1+1+5)// input from AXI bus for additional infor, 8bits messageIbit for TD, lbit for EP, lbit for BCM and 5 bit for typecode, 3bits TC, 2 bits attr,/else
//'define SLV MISC INFO WD(1+ 8 + 3 + 2 +1+1+1+5)// input from AXI bus for additional infor, 8bits message codelbit for BCM and 5 bit for type3bits Tc, 2 bits attr.lbit for TD. lbit for EP.//endif
/////ATOMIC OPERATIONS
////////////////////////////////////////////////define AXI ATOP LOAD LE6'b100o0
------INBOUND BUS DEFINITION-------
---------------------
------
------------------------------
defineINBD HDR PNP RANGE HV LOWINBD HDR PNP RANGE DV LOWdefinedefineINBD HDR PNP RANGE EOT LOWdefineINBD HDR PNP RANGE SEQ LOWdefineINBD HDR PNP RANGE DWEN LOWdefineINBD HDR PNP RANGE DLLP ABORT LOWdefineINBD HDR PNP RANGE TLP ABORT LOWdefineINBD HDR PNP RANGE ECRC ABORT LOWdefineINBD HDR PNP RANGE FMT LOWdefineINBD HDR PNP RANGE TYPE LOW
o
12
3
CC AMBA TLP SEQ WD +3CC AMBA TLP SEO WD +CX NW +3CC AMBA TLP SEO WD +CX NW+4CCAMBATLP SEQ WD+CXNW+5CCAMBA TLP SEQ WD +CXNW+6CC AMBA TLP SEQ WD +CXNW +8CC AMBA TLP SEQ WD +CX NW +13CC AMBA TLP SEO WD +CXNW+1615'ATS RX ENABLE VALUE +CC AMBA TLP SEO WD +CX NW +FLT Q ATTR WIDTH +3*'ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CX NW +FLT Q ATTR WIDTH + 15+CC AMBA TLP SEQ WD +CX NW +FLT Q ATTR WIDTH +163*ATS RX ENABLE VALUE3*ATS RX ENABLE VALUE+CC AMBA TLP SEQ WD +CX NW +FLT Q ATTR WIDTH +323*ATS RX ENABLE VALUE +CC AMBA TLP SEO WD +CX NW +FLT O ATTR WIDTH
defineINBD HDR PNP RANGE TC LOWdefineINBD HDR PNP RANGE ATTR LOWdefineINBD HDR PNP RANGE ATS LOWdefineINBD HDR PNP RANGE NW LOWdefineINBD HDR PNP RANGE REQID LOW
defineINBD HDR PNP RANGE TAG LOWdefineINBD HDR PNP RANGE LOOKUP ID LOW
CX TAGSIZE + 32
define INBD HDR PNP RANGE FUNC NUM LOW3*'ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CX NW +FLT Q ATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD +32define INBD HDR PNP RANGE TD LOW3*ATS RXENABLE VALUE + CC AMBA TLP SEQ WD +CX NFUNC WD +CX NW +FLTQ ATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD +323*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CX NFUNC WD +CX NW +define INBD HDR PNP RANGE POISONED LOWFLT Q ATTR WIDTH +CX TAG SIZE+CX REMOTE MAX TAGS WD+33define INBD HDR PNP RANGE DW LEN LOW3*ATS RX ENABLE VALUE - CC AMBA TLP SEO WD +CX NFUNC WD +CX NW +FLT O ATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD + 34define INBD HDR PNP RANGE FIRST BE LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CX NFUNC WD +CX NW +FLT O ATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD + 44define INBD HDR PNP RANGE LAST BE LOW3*'ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CX NFUNC WD +CX NW +FLT OATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD +483*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CX NFUNC WD +CX NW +define INBD HDR PNP RANGE ADDR LOWFLT Q ATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD + 52define INBD HDR PNP RANGE ROM IN RANGE LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CC CORE ADDR BUS WD +CX NFUNC WD +'CX NW +ELT O ATTR WIDTH +CX TAG SIZE +CX REMOTE MAX TAGS WD + 52define INBD HDR PNP RANGE IOREQ IN RANGE LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CC CORE ADDR BUS WD +CX NFUNC WD + 'CX NW +FLT O ATTR WIDTH + CX TAG SIZE -CX REMOTE MAX AGS WD + 53define INBD HDR PNP RANGE IN MEMBAR RANGE LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEO WD +CC CORE ADDR BUS WD +CX NFUNC WD +'CX NW +FLT Q ATTR WIDTH + CX TAG SIZE +CX REMOTE MAX TAGS WD + 543*ATS RX ENABLE VALUE +CC AMBA TLP SEO WD +CC CORE ADDR BUS WD +define INBD HDR PNP RANGE TPH SET LOWCX NFUNC WD + 'CX NW + CX TPH ENABLE VALUE + FLT O ATTR WIDTH + CX TAG SIZE + CX REMOTE MAX TAGS WD + 56define INBD HDR PNP RANGE TPH PH LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEO WD +CC CORE ADDR BUS WD+CX NFUNC WD + 'CX NW + 9*'CX TPH ENABLE VALUE + FLT O ATTR WIDTH + CX TAG SIZE + CX REMOTE MAX TAS WD + 56define INBD HDR PNP RANGE TPH TH LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CC CORE ADDR BUS WD +CX NFUNC WD + 'CX NW + 11'CX TPH ENABLE VALUE + FLT O ATTR WIDTH - CX TAG SIZE + CX REMOTE MAX TAGS WD + 56define INBD HDR PNP RANGE MEM TYPE LOW3ATS RX ENABLE VALUE +CC AMBA TLP SEO WD +CC CORE ADDR BUS WD+CX NFUNC WD + 'CX NW + 11'CX TPH ENABLE VALUE + FLT  ATTR WIDTH + CX TAG SIZE + CX REMOTE MAX TAGS WD + 573*ATS RX ENABLE VALUE +CC AMBA TLP SEQ WD +CC CORE ADDR BUS WD +define INBD HDR PNP RANGE VC NUM LOWCX NFUNC WD + 'CX MM + 11'CX TPH ENABLE VALUE + RADN SEG BUF VALUE*'DC MULTI NC VALUE - FLT O ATTR VTDTH - CX TAG STZE +CXREMOTE MAX TAGS WD + 57define INBD HDR PNP RANGE BCM LOW3*ATS RX ENABLE VALUE +CC AMBA TLP SEO WD -CC CORE ADDR BUS WD +CX NFUNC WD + 'CX NW + 11'CX TPH ENABLE VALUE + RADM SEG BUF VALUEDC MULTI VC VALUEI'CX NVC LOG2  1)+RADM SEG BUF VALUE*'DC MULTI VC VALUE + FLT O ATTR WIDTH + RADM SEG BUF VALUE + CX TAG SIZE + CX REMOTE MAX TAGS WD + 57
////I/1// PCIe ATS Translation Response message fieldsdefine DC PCIE ATS TRSP TADDR WD 52
II/I///////////
////////////
/ ATS Invalidate Completion Message Fields
//////////////////////////////////////////////I/I////////////define DC PCIE ATS INV COMP ITAG VEC MSB 31define DC PCIE ATS INV COMP ITAG VEC WD 32
define DC PCIE ATS INV COMP CC MSB 34
define DC PCIE ATS INV COMP CC WD 3
////////////////////////////////////////////I///////////// PCIe Page Response messagedefine DC PCIE ATS PRSP RESP CODE WD 4
/ RESP CODE field encodingdefine DC PCIE PCOMP RSPCODE SUCCESS 4'b0000
define DC PCIE PCOMP RSPCODE INV REQ 4'b0001define DC PCIE PCOMP RSPCODE FAIL 4'b1111
/////////////////////////////////////////
//DTIM Register Fields
define DC DTIM ROOT PORT ID WD 16
define DC DTIM TOK TRANS REQ WD 8
define DC DTIM IREQ TO RNG WD 3
define DC DTIM FLUSH IREQ SID WD 16
define DC DTIM CONDIS REQ WD 2
/ AXI4-Stream Master Message priority, lowest value has highest priority
define DC DTIM SM PRIOR WEIGHT WD 3
define DC TRANS REO MSG PRIORITY 3 b100
define DC PAGE REQ MSG PRIORITY 3'b010
define DC SYNC ACK MSG PRIORITY 3'b001define DC INV ACK MSG PRIORITY 3'b000
define DC DTIM TREQ QOS WD 4
define DC DTIM MSI ADDR UPR WD 32
define DC DTIM MSI ADDR LWR WD 30
define DC DTIM MSI DATA WD 32
define DC DTIM ERR IREQ OPCODE WD 8
define DC DTIM ERR IREQ TO ITAG WD 5
define DC DTIM ERR IREQ TO SID LWR WD 16
define DC DTIM ERR ICPL UC ITAG WD 5
define DC DTIM ERR ICPL UC REQ ID WD 16
define DC DTIM ERR TRESP UR TID WD 8
define DC DTIM TOK TREQ GNT WD 8
define DC DTIM OAS WD 4
define DC DTIM CONDIS STATE WD 2
define DC DTIM IREQ TMR TO WD 16define DC DTIM IREQ TMR TO SF WD 2
endif1/
GUARD AMBA DEFS SVH